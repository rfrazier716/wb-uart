`default_nettype none //flags an error if you haven't defined a wire


// A basic uart example that transmits a message every second

module hello_uart(
    input wire i_clk, // The system clock
    output wire o_tx_w, // uart TX wire
    output wire i_rx_w // uart Tx wire
);



endmodule;